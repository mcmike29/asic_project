VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dynamic_noise_reduction
  CLASS BLOCK ;
  FOREIGN dynamic_noise_reduction ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 507.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 -9.470 514.390 -6.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 504.130 514.390 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 511.290 -9.470 514.390 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.570 -9.470 30.670 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 127.570 -9.470 130.670 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 227.570 -9.470 230.670 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 327.570 -9.470 330.670 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 427.570 -9.470 430.670 507.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 32.930 514.390 36.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 132.930 514.390 136.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 232.930 514.390 236.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 332.930 514.390 336.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 432.930 514.390 436.030 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 502.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 -4.670 509.590 -1.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 499.330 509.590 502.430 ;
    END
    PORT
      LAYER met4 ;
        RECT 506.490 -4.670 509.590 502.430 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 -9.470 12.070 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.970 -9.470 112.070 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.970 -9.470 212.070 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.970 -9.470 312.070 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.970 -9.470 412.070 507.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 14.330 514.390 17.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 114.330 514.390 117.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 214.330 514.390 217.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 314.330 514.390 317.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 414.330 514.390 417.430 ;
    END
  END VPWR
  PIN alpha[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 102.040 500.000 102.640 ;
    END
  END alpha[0]
  PIN alpha[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END alpha[10]
  PIN alpha[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END alpha[11]
  PIN alpha[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END alpha[12]
  PIN alpha[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END alpha[13]
  PIN alpha[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END alpha[14]
  PIN alpha[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END alpha[15]
  PIN alpha[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 105.440 500.000 106.040 ;
    END
  END alpha[1]
  PIN alpha[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 108.840 500.000 109.440 ;
    END
  END alpha[2]
  PIN alpha[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 88.440 500.000 89.040 ;
    END
  END alpha[3]
  PIN alpha[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 91.840 500.000 92.440 ;
    END
  END alpha[4]
  PIN alpha[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 95.240 500.000 95.840 ;
    END
  END alpha[5]
  PIN alpha[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END alpha[6]
  PIN alpha[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END alpha[7]
  PIN alpha[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END alpha[8]
  PIN alpha[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END alpha[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END reset
  PIN x_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 217.640 500.000 218.240 ;
    END
  END x_in[0]
  PIN x_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END x_in[10]
  PIN x_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END x_in[11]
  PIN x_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END x_in[12]
  PIN x_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END x_in[13]
  PIN x_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END x_in[14]
  PIN x_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END x_in[15]
  PIN x_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 214.240 500.000 214.840 ;
    END
  END x_in[1]
  PIN x_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 204.040 500.000 204.640 ;
    END
  END x_in[2]
  PIN x_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 187.040 500.000 187.640 ;
    END
  END x_in[3]
  PIN x_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 180.240 500.000 180.840 ;
    END
  END x_in[4]
  PIN x_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 163.240 500.000 163.840 ;
    END
  END x_in[5]
  PIN x_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 156.440 500.000 157.040 ;
    END
  END x_in[6]
  PIN x_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END x_in[7]
  PIN x_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END x_in[8]
  PIN x_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END x_in[9]
  PIN y_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 255.040 500.000 255.640 ;
    END
  END y_out[0]
  PIN y_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END y_out[10]
  PIN y_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END y_out[11]
  PIN y_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 289.890 496.000 290.170 500.000 ;
    END
  END y_out[12]
  PIN y_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END y_out[13]
  PIN y_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END y_out[14]
  PIN y_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END y_out[15]
  PIN y_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 221.040 500.000 221.640 ;
    END
  END y_out[1]
  PIN y_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 268.640 500.000 269.240 ;
    END
  END y_out[2]
  PIN y_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 272.040 500.000 272.640 ;
    END
  END y_out[3]
  PIN y_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 275.440 500.000 276.040 ;
    END
  END y_out[4]
  PIN y_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 234.640 500.000 235.240 ;
    END
  END y_out[5]
  PIN y_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 224.440 500.000 225.040 ;
    END
  END y_out[6]
  PIN y_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 402.590 496.000 402.870 500.000 ;
    END
  END y_out[7]
  PIN y_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 380.050 496.000 380.330 500.000 ;
    END
  END y_out[8]
  PIN y_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 376.830 496.000 377.110 500.000 ;
    END
  END y_out[9]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 494.230 487.070 ;
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 0.530 10.640 494.040 487.120 ;
      LAYER met2 ;
        RECT 0.550 495.720 289.610 496.810 ;
        RECT 290.450 495.720 376.550 496.810 ;
        RECT 377.390 495.720 379.770 496.810 ;
        RECT 380.610 495.720 402.310 496.810 ;
        RECT 403.150 495.720 492.570 496.810 ;
        RECT 0.550 4.280 492.570 495.720 ;
        RECT 0.550 4.000 70.650 4.280 ;
        RECT 71.490 4.000 73.870 4.280 ;
        RECT 74.710 4.000 77.090 4.280 ;
        RECT 77.930 4.000 80.310 4.280 ;
        RECT 81.150 4.000 83.530 4.280 ;
        RECT 84.370 4.000 99.630 4.280 ;
        RECT 100.470 4.000 118.950 4.280 ;
        RECT 119.790 4.000 122.170 4.280 ;
        RECT 123.010 4.000 135.050 4.280 ;
        RECT 135.890 4.000 138.270 4.280 ;
        RECT 139.110 4.000 144.710 4.280 ;
        RECT 145.550 4.000 167.250 4.280 ;
        RECT 168.090 4.000 492.570 4.280 ;
      LAYER met3 ;
        RECT 0.525 419.240 496.000 487.045 ;
        RECT 4.400 417.840 496.000 419.240 ;
        RECT 0.525 415.840 496.000 417.840 ;
        RECT 4.400 414.440 496.000 415.840 ;
        RECT 0.525 405.640 496.000 414.440 ;
        RECT 4.400 404.240 496.000 405.640 ;
        RECT 0.525 392.040 496.000 404.240 ;
        RECT 4.400 390.640 496.000 392.040 ;
        RECT 0.525 388.640 496.000 390.640 ;
        RECT 4.400 387.240 496.000 388.640 ;
        RECT 0.525 378.440 496.000 387.240 ;
        RECT 4.400 377.040 496.000 378.440 ;
        RECT 0.525 375.040 496.000 377.040 ;
        RECT 4.400 373.640 496.000 375.040 ;
        RECT 0.525 364.840 496.000 373.640 ;
        RECT 4.400 363.440 496.000 364.840 ;
        RECT 0.525 344.440 496.000 363.440 ;
        RECT 4.400 343.040 496.000 344.440 ;
        RECT 0.525 330.840 496.000 343.040 ;
        RECT 4.400 329.440 496.000 330.840 ;
        RECT 0.525 307.040 496.000 329.440 ;
        RECT 4.400 305.640 496.000 307.040 ;
        RECT 0.525 293.440 496.000 305.640 ;
        RECT 4.400 292.040 496.000 293.440 ;
        RECT 0.525 283.240 496.000 292.040 ;
        RECT 4.400 281.840 496.000 283.240 ;
        RECT 0.525 276.440 496.000 281.840 ;
        RECT 0.525 275.040 495.600 276.440 ;
        RECT 0.525 273.040 496.000 275.040 ;
        RECT 4.400 271.640 495.600 273.040 ;
        RECT 0.525 269.640 496.000 271.640 ;
        RECT 0.525 268.240 495.600 269.640 ;
        RECT 0.525 256.040 496.000 268.240 ;
        RECT 0.525 254.640 495.600 256.040 ;
        RECT 0.525 235.640 496.000 254.640 ;
        RECT 0.525 234.240 495.600 235.640 ;
        RECT 0.525 225.440 496.000 234.240 ;
        RECT 0.525 224.040 495.600 225.440 ;
        RECT 0.525 222.040 496.000 224.040 ;
        RECT 0.525 220.640 495.600 222.040 ;
        RECT 0.525 218.640 496.000 220.640 ;
        RECT 0.525 217.240 495.600 218.640 ;
        RECT 0.525 215.240 496.000 217.240 ;
        RECT 0.525 213.840 495.600 215.240 ;
        RECT 0.525 205.040 496.000 213.840 ;
        RECT 0.525 203.640 495.600 205.040 ;
        RECT 0.525 188.040 496.000 203.640 ;
        RECT 0.525 186.640 495.600 188.040 ;
        RECT 0.525 181.240 496.000 186.640 ;
        RECT 0.525 179.840 495.600 181.240 ;
        RECT 0.525 164.240 496.000 179.840 ;
        RECT 0.525 162.840 495.600 164.240 ;
        RECT 0.525 157.440 496.000 162.840 ;
        RECT 0.525 156.040 495.600 157.440 ;
        RECT 0.525 109.840 496.000 156.040 ;
        RECT 0.525 108.440 495.600 109.840 ;
        RECT 0.525 106.440 496.000 108.440 ;
        RECT 0.525 105.040 495.600 106.440 ;
        RECT 0.525 103.040 496.000 105.040 ;
        RECT 0.525 101.640 495.600 103.040 ;
        RECT 0.525 96.240 496.000 101.640 ;
        RECT 0.525 94.840 495.600 96.240 ;
        RECT 0.525 92.840 496.000 94.840 ;
        RECT 0.525 91.440 495.600 92.840 ;
        RECT 0.525 89.440 496.000 91.440 ;
        RECT 0.525 88.040 495.600 89.440 ;
        RECT 0.525 10.715 496.000 88.040 ;
      LAYER met4 ;
        RECT 142.895 107.615 208.570 332.345 ;
        RECT 212.470 107.615 227.170 332.345 ;
        RECT 231.070 107.615 308.570 332.345 ;
        RECT 312.470 107.615 327.170 332.345 ;
        RECT 331.070 107.615 408.570 332.345 ;
        RECT 412.470 107.615 413.705 332.345 ;
  END
END dynamic_noise_reduction
END LIBRARY

