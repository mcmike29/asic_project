VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dynamic_noise_reduction
  CLASS BLOCK ;
  FOREIGN dynamic_noise_reduction ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 1000.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 1007.710 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 -9.470 1014.410 -6.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1004.610 1014.410 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 1011.310 -9.470 1014.410 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.570 -9.470 30.670 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 127.570 -9.470 130.670 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 227.570 -9.470 230.670 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 327.570 -9.470 330.670 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 427.570 -9.470 430.670 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 527.570 -9.470 530.670 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 627.570 -9.470 630.670 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 727.570 -9.470 730.670 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 827.570 -9.470 830.670 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.570 -9.470 930.670 1007.710 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 32.930 1014.410 36.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 132.930 1014.410 136.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 232.930 1014.410 236.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 332.930 1014.410 336.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 432.930 1014.410 436.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 532.930 1014.410 536.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 632.930 1014.410 636.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 732.930 1014.410 736.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 832.930 1014.410 836.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 932.930 1014.410 936.030 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 1002.910 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 -4.670 1009.610 -1.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 999.810 1009.610 1002.910 ;
    END
    PORT
      LAYER met4 ;
        RECT 1006.510 -4.670 1009.610 1002.910 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 -9.470 12.070 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.970 -9.470 112.070 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.970 -9.470 212.070 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.970 -9.470 312.070 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.970 -9.470 412.070 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.970 -9.470 512.070 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 608.970 -9.470 612.070 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 708.970 -9.470 712.070 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 808.970 -9.470 812.070 1007.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 -9.470 912.070 1007.710 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 14.330 1014.410 17.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 114.330 1014.410 117.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 214.330 1014.410 217.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 314.330 1014.410 317.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 414.330 1014.410 417.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 514.330 1014.410 517.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 614.330 1014.410 617.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 714.330 1014.410 717.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 814.330 1014.410 817.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 914.330 1014.410 917.430 ;
    END
  END VPWR
  PIN alpha[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 333.240 1000.000 333.840 ;
    END
  END alpha[0]
  PIN alpha[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END alpha[10]
  PIN alpha[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END alpha[11]
  PIN alpha[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END alpha[12]
  PIN alpha[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END alpha[13]
  PIN alpha[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END alpha[14]
  PIN alpha[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END alpha[15]
  PIN alpha[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 336.640 1000.000 337.240 ;
    END
  END alpha[1]
  PIN alpha[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 340.040 1000.000 340.640 ;
    END
  END alpha[2]
  PIN alpha[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 343.440 1000.000 344.040 ;
    END
  END alpha[3]
  PIN alpha[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 346.840 1000.000 347.440 ;
    END
  END alpha[4]
  PIN alpha[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 350.240 1000.000 350.840 ;
    END
  END alpha[5]
  PIN alpha[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 329.840 1000.000 330.440 ;
    END
  END alpha[6]
  PIN alpha[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 353.640 1000.000 354.240 ;
    END
  END alpha[7]
  PIN alpha[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END alpha[8]
  PIN alpha[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END alpha[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END reset
  PIN x_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 448.840 1000.000 449.440 ;
    END
  END x_in[0]
  PIN x_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END x_in[10]
  PIN x_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END x_in[11]
  PIN x_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END x_in[12]
  PIN x_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END x_in[13]
  PIN x_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END x_in[14]
  PIN x_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END x_in[15]
  PIN x_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 438.640 1000.000 439.240 ;
    END
  END x_in[1]
  PIN x_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 431.840 1000.000 432.440 ;
    END
  END x_in[2]
  PIN x_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 425.040 1000.000 425.640 ;
    END
  END x_in[3]
  PIN x_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 408.040 1000.000 408.640 ;
    END
  END x_in[4]
  PIN x_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 397.840 1000.000 398.440 ;
    END
  END x_in[5]
  PIN x_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 384.240 1000.000 384.840 ;
    END
  END x_in[6]
  PIN x_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 374.040 1000.000 374.640 ;
    END
  END x_in[7]
  PIN x_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 367.240 1000.000 367.840 ;
    END
  END x_in[8]
  PIN x_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 357.040 1000.000 357.640 ;
    END
  END x_in[9]
  PIN y_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 496.440 1000.000 497.040 ;
    END
  END y_out[0]
  PIN y_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END y_out[10]
  PIN y_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END y_out[11]
  PIN y_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END y_out[12]
  PIN y_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END y_out[13]
  PIN y_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END y_out[14]
  PIN y_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END y_out[15]
  PIN y_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 462.440 1000.000 463.040 ;
    END
  END y_out[1]
  PIN y_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 785.770 996.000 786.050 1000.000 ;
    END
  END y_out[2]
  PIN y_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 782.550 996.000 782.830 1000.000 ;
    END
  END y_out[3]
  PIN y_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 779.330 996.000 779.610 1000.000 ;
    END
  END y_out[4]
  PIN y_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 753.570 996.000 753.850 1000.000 ;
    END
  END y_out[5]
  PIN y_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 750.350 996.000 750.630 1000.000 ;
    END
  END y_out[6]
  PIN y_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 705.270 996.000 705.550 1000.000 ;
    END
  END y_out[7]
  PIN y_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END y_out[8]
  PIN y_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END y_out[9]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 994.250 987.550 ;
      LAYER li1 ;
        RECT 5.520 10.795 994.060 987.445 ;
      LAYER met1 ;
        RECT 0.530 10.640 994.060 987.600 ;
      LAYER met2 ;
        RECT 0.550 995.720 704.990 996.610 ;
        RECT 705.830 995.720 750.070 996.610 ;
        RECT 750.910 995.720 753.290 996.610 ;
        RECT 754.130 995.720 779.050 996.610 ;
        RECT 779.890 995.720 782.270 996.610 ;
        RECT 783.110 995.720 785.490 996.610 ;
        RECT 786.330 995.720 992.590 996.610 ;
        RECT 0.550 4.280 992.590 995.720 ;
        RECT 0.550 4.000 189.790 4.280 ;
        RECT 190.630 4.000 193.010 4.280 ;
        RECT 193.850 4.000 196.230 4.280 ;
        RECT 197.070 4.000 199.450 4.280 ;
        RECT 200.290 4.000 212.330 4.280 ;
        RECT 213.170 4.000 241.310 4.280 ;
        RECT 242.150 4.000 263.850 4.280 ;
        RECT 264.690 4.000 992.590 4.280 ;
      LAYER met3 ;
        RECT 0.525 684.440 996.000 987.525 ;
        RECT 4.400 683.040 996.000 684.440 ;
        RECT 0.525 681.040 996.000 683.040 ;
        RECT 4.400 679.640 996.000 681.040 ;
        RECT 0.525 677.640 996.000 679.640 ;
        RECT 4.400 676.240 996.000 677.640 ;
        RECT 0.525 674.240 996.000 676.240 ;
        RECT 4.400 672.840 996.000 674.240 ;
        RECT 0.525 670.840 996.000 672.840 ;
        RECT 4.400 669.440 996.000 670.840 ;
        RECT 0.525 667.440 996.000 669.440 ;
        RECT 4.400 666.040 996.000 667.440 ;
        RECT 0.525 664.040 996.000 666.040 ;
        RECT 4.400 662.640 996.000 664.040 ;
        RECT 0.525 660.640 996.000 662.640 ;
        RECT 4.400 659.240 996.000 660.640 ;
        RECT 0.525 657.240 996.000 659.240 ;
        RECT 4.400 655.840 996.000 657.240 ;
        RECT 0.525 650.440 996.000 655.840 ;
        RECT 4.400 649.040 996.000 650.440 ;
        RECT 0.525 647.040 996.000 649.040 ;
        RECT 4.400 645.640 996.000 647.040 ;
        RECT 0.525 643.640 996.000 645.640 ;
        RECT 4.400 642.240 996.000 643.640 ;
        RECT 0.525 589.240 996.000 642.240 ;
        RECT 4.400 587.840 996.000 589.240 ;
        RECT 0.525 555.240 996.000 587.840 ;
        RECT 4.400 553.840 996.000 555.240 ;
        RECT 0.525 538.240 996.000 553.840 ;
        RECT 4.400 536.840 996.000 538.240 ;
        RECT 0.525 524.640 996.000 536.840 ;
        RECT 4.400 523.240 996.000 524.640 ;
        RECT 0.525 507.640 996.000 523.240 ;
        RECT 4.400 506.240 996.000 507.640 ;
        RECT 0.525 497.440 996.000 506.240 ;
        RECT 0.525 496.040 995.600 497.440 ;
        RECT 0.525 463.440 996.000 496.040 ;
        RECT 0.525 462.040 995.600 463.440 ;
        RECT 0.525 449.840 996.000 462.040 ;
        RECT 0.525 448.440 995.600 449.840 ;
        RECT 0.525 439.640 996.000 448.440 ;
        RECT 0.525 438.240 995.600 439.640 ;
        RECT 0.525 432.840 996.000 438.240 ;
        RECT 0.525 431.440 995.600 432.840 ;
        RECT 0.525 426.040 996.000 431.440 ;
        RECT 0.525 424.640 995.600 426.040 ;
        RECT 0.525 409.040 996.000 424.640 ;
        RECT 0.525 407.640 995.600 409.040 ;
        RECT 0.525 398.840 996.000 407.640 ;
        RECT 0.525 397.440 995.600 398.840 ;
        RECT 0.525 385.240 996.000 397.440 ;
        RECT 0.525 383.840 995.600 385.240 ;
        RECT 0.525 375.040 996.000 383.840 ;
        RECT 0.525 373.640 995.600 375.040 ;
        RECT 0.525 368.240 996.000 373.640 ;
        RECT 0.525 366.840 995.600 368.240 ;
        RECT 0.525 358.040 996.000 366.840 ;
        RECT 0.525 356.640 995.600 358.040 ;
        RECT 0.525 354.640 996.000 356.640 ;
        RECT 0.525 353.240 995.600 354.640 ;
        RECT 0.525 351.240 996.000 353.240 ;
        RECT 0.525 349.840 995.600 351.240 ;
        RECT 0.525 347.840 996.000 349.840 ;
        RECT 0.525 346.440 995.600 347.840 ;
        RECT 0.525 344.440 996.000 346.440 ;
        RECT 0.525 343.040 995.600 344.440 ;
        RECT 0.525 341.040 996.000 343.040 ;
        RECT 0.525 339.640 995.600 341.040 ;
        RECT 0.525 337.640 996.000 339.640 ;
        RECT 0.525 336.240 995.600 337.640 ;
        RECT 0.525 334.240 996.000 336.240 ;
        RECT 0.525 332.840 995.600 334.240 ;
        RECT 0.525 330.840 996.000 332.840 ;
        RECT 0.525 329.440 995.600 330.840 ;
        RECT 0.525 10.715 996.000 329.440 ;
      LAYER met4 ;
        RECT 3.975 357.855 8.570 678.465 ;
        RECT 12.470 357.855 27.170 678.465 ;
        RECT 31.070 357.855 108.570 678.465 ;
        RECT 112.470 357.855 127.170 678.465 ;
        RECT 131.070 357.855 208.570 678.465 ;
        RECT 212.470 357.855 227.170 678.465 ;
        RECT 231.070 357.855 308.570 678.465 ;
        RECT 312.470 357.855 327.170 678.465 ;
        RECT 331.070 357.855 408.570 678.465 ;
        RECT 412.470 357.855 427.170 678.465 ;
        RECT 431.070 357.855 508.570 678.465 ;
        RECT 512.470 357.855 527.170 678.465 ;
        RECT 531.070 357.855 608.570 678.465 ;
        RECT 612.470 357.855 627.170 678.465 ;
        RECT 631.070 357.855 708.570 678.465 ;
        RECT 712.470 357.855 727.170 678.465 ;
        RECT 731.070 357.855 808.570 678.465 ;
        RECT 812.470 357.855 827.170 678.465 ;
        RECT 831.070 357.855 908.570 678.465 ;
        RECT 912.470 357.855 927.170 678.465 ;
        RECT 931.070 357.855 982.265 678.465 ;
  END
END dynamic_noise_reduction
END LIBRARY

