VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dynamic_noise_reduction
  CLASS BLOCK ;
  FOREIGN dynamic_noise_reduction ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 507.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 -9.470 514.390 -6.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 504.130 514.390 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 511.290 -9.470 514.390 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.570 -9.470 30.670 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 127.570 -9.470 130.670 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 227.570 -9.470 230.670 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 327.570 -9.470 330.670 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 427.570 -9.470 430.670 507.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 32.930 514.390 36.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 132.930 514.390 136.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 232.930 514.390 236.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 332.930 514.390 336.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 432.930 514.390 436.030 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 502.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 -4.670 509.590 -1.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 499.330 509.590 502.430 ;
    END
    PORT
      LAYER met4 ;
        RECT 506.490 -4.670 509.590 502.430 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 -9.470 12.070 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.970 -9.470 112.070 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.970 -9.470 212.070 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.970 -9.470 312.070 507.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.970 -9.470 412.070 507.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 14.330 514.390 17.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 114.330 514.390 117.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 214.330 514.390 217.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 314.330 514.390 317.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 414.330 514.390 417.430 ;
    END
  END VPWR
  PIN alpha[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 88.440 500.000 89.040 ;
    END
  END alpha[0]
  PIN alpha[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END alpha[10]
  PIN alpha[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END alpha[11]
  PIN alpha[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END alpha[12]
  PIN alpha[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END alpha[13]
  PIN alpha[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END alpha[14]
  PIN alpha[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END alpha[15]
  PIN alpha[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 91.840 500.000 92.440 ;
    END
  END alpha[1]
  PIN alpha[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 95.240 500.000 95.840 ;
    END
  END alpha[2]
  PIN alpha[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 98.640 500.000 99.240 ;
    END
  END alpha[3]
  PIN alpha[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 102.040 500.000 102.640 ;
    END
  END alpha[4]
  PIN alpha[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 105.440 500.000 106.040 ;
    END
  END alpha[5]
  PIN alpha[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 85.040 500.000 85.640 ;
    END
  END alpha[6]
  PIN alpha[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END alpha[7]
  PIN alpha[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END alpha[8]
  PIN alpha[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END alpha[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END reset
  PIN x_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 210.840 500.000 211.440 ;
    END
  END x_in[0]
  PIN x_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END x_in[10]
  PIN x_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END x_in[11]
  PIN x_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END x_in[12]
  PIN x_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END x_in[13]
  PIN x_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END x_in[14]
  PIN x_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END x_in[15]
  PIN x_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 200.640 500.000 201.240 ;
    END
  END x_in[1]
  PIN x_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 187.040 500.000 187.640 ;
    END
  END x_in[2]
  PIN x_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 180.240 500.000 180.840 ;
    END
  END x_in[3]
  PIN x_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 170.040 500.000 170.640 ;
    END
  END x_in[4]
  PIN x_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 159.840 500.000 160.440 ;
    END
  END x_in[5]
  PIN x_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 149.640 500.000 150.240 ;
    END
  END x_in[6]
  PIN x_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END x_in[7]
  PIN x_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END x_in[8]
  PIN x_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END x_in[9]
  PIN y_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 251.640 500.000 252.240 ;
    END
  END y_out[0]
  PIN y_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 228.710 496.000 228.990 500.000 ;
    END
  END y_out[10]
  PIN y_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END y_out[11]
  PIN y_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END y_out[12]
  PIN y_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END y_out[13]
  PIN y_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END y_out[14]
  PIN y_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END y_out[15]
  PIN y_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 227.840 500.000 228.440 ;
    END
  END y_out[1]
  PIN y_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 244.840 500.000 245.440 ;
    END
  END y_out[2]
  PIN y_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 255.040 500.000 255.640 ;
    END
  END y_out[3]
  PIN y_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 258.440 500.000 259.040 ;
    END
  END y_out[4]
  PIN y_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 241.440 500.000 242.040 ;
    END
  END y_out[5]
  PIN y_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 224.440 500.000 225.040 ;
    END
  END y_out[6]
  PIN y_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 193.840 500.000 194.440 ;
    END
  END y_out[7]
  PIN y_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 386.490 496.000 386.770 500.000 ;
    END
  END y_out[8]
  PIN y_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 370.390 496.000 370.670 500.000 ;
    END
  END y_out[9]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 494.230 487.070 ;
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 0.530 10.640 494.040 487.120 ;
      LAYER met2 ;
        RECT 0.550 495.720 228.430 496.810 ;
        RECT 229.270 495.720 370.110 496.810 ;
        RECT 370.950 495.720 386.210 496.810 ;
        RECT 387.050 495.720 492.570 496.810 ;
        RECT 0.550 4.280 492.570 495.720 ;
        RECT 0.550 4.000 48.110 4.280 ;
        RECT 48.950 4.000 51.330 4.280 ;
        RECT 52.170 4.000 54.550 4.280 ;
        RECT 55.390 4.000 57.770 4.280 ;
        RECT 58.610 4.000 80.310 4.280 ;
        RECT 81.150 4.000 96.410 4.280 ;
        RECT 97.250 4.000 115.730 4.280 ;
        RECT 116.570 4.000 118.950 4.280 ;
        RECT 119.790 4.000 125.390 4.280 ;
        RECT 126.230 4.000 131.830 4.280 ;
        RECT 132.670 4.000 170.470 4.280 ;
        RECT 171.310 4.000 492.570 4.280 ;
      LAYER met3 ;
        RECT 0.525 405.640 496.000 487.045 ;
        RECT 4.400 404.240 496.000 405.640 ;
        RECT 0.525 398.840 496.000 404.240 ;
        RECT 4.400 397.440 496.000 398.840 ;
        RECT 0.525 395.440 496.000 397.440 ;
        RECT 4.400 394.040 496.000 395.440 ;
        RECT 0.525 392.040 496.000 394.040 ;
        RECT 4.400 390.640 496.000 392.040 ;
        RECT 0.525 378.440 496.000 390.640 ;
        RECT 4.400 377.040 496.000 378.440 ;
        RECT 0.525 371.640 496.000 377.040 ;
        RECT 4.400 370.240 496.000 371.640 ;
        RECT 0.525 368.240 496.000 370.240 ;
        RECT 4.400 366.840 496.000 368.240 ;
        RECT 0.525 354.640 496.000 366.840 ;
        RECT 4.400 353.240 496.000 354.640 ;
        RECT 0.525 351.240 496.000 353.240 ;
        RECT 4.400 349.840 496.000 351.240 ;
        RECT 0.525 344.440 496.000 349.840 ;
        RECT 4.400 343.040 496.000 344.440 ;
        RECT 0.525 293.440 496.000 343.040 ;
        RECT 4.400 292.040 496.000 293.440 ;
        RECT 0.525 269.640 496.000 292.040 ;
        RECT 4.400 268.240 496.000 269.640 ;
        RECT 0.525 259.440 496.000 268.240 ;
        RECT 4.400 258.040 495.600 259.440 ;
        RECT 0.525 256.040 496.000 258.040 ;
        RECT 4.400 254.640 495.600 256.040 ;
        RECT 0.525 252.640 496.000 254.640 ;
        RECT 0.525 251.240 495.600 252.640 ;
        RECT 0.525 245.840 496.000 251.240 ;
        RECT 0.525 244.440 495.600 245.840 ;
        RECT 0.525 242.440 496.000 244.440 ;
        RECT 0.525 241.040 495.600 242.440 ;
        RECT 0.525 228.840 496.000 241.040 ;
        RECT 0.525 227.440 495.600 228.840 ;
        RECT 0.525 225.440 496.000 227.440 ;
        RECT 0.525 224.040 495.600 225.440 ;
        RECT 0.525 211.840 496.000 224.040 ;
        RECT 0.525 210.440 495.600 211.840 ;
        RECT 0.525 201.640 496.000 210.440 ;
        RECT 0.525 200.240 495.600 201.640 ;
        RECT 0.525 194.840 496.000 200.240 ;
        RECT 0.525 193.440 495.600 194.840 ;
        RECT 0.525 188.040 496.000 193.440 ;
        RECT 0.525 186.640 495.600 188.040 ;
        RECT 0.525 181.240 496.000 186.640 ;
        RECT 0.525 179.840 495.600 181.240 ;
        RECT 0.525 171.040 496.000 179.840 ;
        RECT 0.525 169.640 495.600 171.040 ;
        RECT 0.525 160.840 496.000 169.640 ;
        RECT 0.525 159.440 495.600 160.840 ;
        RECT 0.525 150.640 496.000 159.440 ;
        RECT 0.525 149.240 495.600 150.640 ;
        RECT 0.525 106.440 496.000 149.240 ;
        RECT 0.525 105.040 495.600 106.440 ;
        RECT 0.525 103.040 496.000 105.040 ;
        RECT 0.525 101.640 495.600 103.040 ;
        RECT 0.525 99.640 496.000 101.640 ;
        RECT 0.525 98.240 495.600 99.640 ;
        RECT 0.525 96.240 496.000 98.240 ;
        RECT 0.525 94.840 495.600 96.240 ;
        RECT 0.525 92.840 496.000 94.840 ;
        RECT 0.525 91.440 495.600 92.840 ;
        RECT 0.525 89.440 496.000 91.440 ;
        RECT 0.525 88.040 495.600 89.440 ;
        RECT 0.525 86.040 496.000 88.040 ;
        RECT 0.525 84.640 495.600 86.040 ;
        RECT 0.525 10.715 496.000 84.640 ;
      LAYER met4 ;
        RECT 343.455 155.895 408.570 346.625 ;
        RECT 412.470 155.895 427.170 346.625 ;
        RECT 431.070 155.895 489.145 346.625 ;
  END
END dynamic_noise_reduction
END LIBRARY

